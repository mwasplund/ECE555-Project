library verilog;
use verilog.vl_types.all;
entity \NAND\ is
    port(
        \OUT\           : out    vl_logic;
        IN1             : in     vl_logic;
        IN2             : in     vl_logic
    );
end \NAND\;
