library verilog;
use verilog.vl_types.all;
entity Buffer_1bit is
    port(
        \OUT\           : out    vl_logic;
        \IN\            : in     vl_logic
    );
end Buffer_1bit;
