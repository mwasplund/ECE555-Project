library verilog;
use verilog.vl_types.all;
entity Adder_32bit_nlogic is
    port(
        Cout            : out    vl_logic;
        S0              : out    vl_logic;
        S1              : out    vl_logic;
        S2              : out    vl_logic;
        S3              : out    vl_logic;
        S4              : out    vl_logic;
        S5              : out    vl_logic;
        S6              : out    vl_logic;
        S7              : out    vl_logic;
        S8              : out    vl_logic;
        S9              : out    vl_logic;
        S10             : out    vl_logic;
        S11             : out    vl_logic;
        S12             : out    vl_logic;
        S13             : out    vl_logic;
        S14             : out    vl_logic;
        S15             : out    vl_logic;
        S16             : out    vl_logic;
        S17             : out    vl_logic;
        S18             : out    vl_logic;
        S19             : out    vl_logic;
        S20             : out    vl_logic;
        S21             : out    vl_logic;
        S22             : out    vl_logic;
        S23             : out    vl_logic;
        S24             : out    vl_logic;
        S25             : out    vl_logic;
        S26             : out    vl_logic;
        S27             : out    vl_logic;
        S28             : out    vl_logic;
        S29             : out    vl_logic;
        S30             : out    vl_logic;
        S31             : out    vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        A4              : in     vl_logic;
        A5              : in     vl_logic;
        A6              : in     vl_logic;
        A7              : in     vl_logic;
        A8              : in     vl_logic;
        A9              : in     vl_logic;
        A10             : in     vl_logic;
        A11             : in     vl_logic;
        A12             : in     vl_logic;
        A13             : in     vl_logic;
        A14             : in     vl_logic;
        A15             : in     vl_logic;
        A16             : in     vl_logic;
        A17             : in     vl_logic;
        A18             : in     vl_logic;
        A19             : in     vl_logic;
        A20             : in     vl_logic;
        A21             : in     vl_logic;
        A22             : in     vl_logic;
        A23             : in     vl_logic;
        A24             : in     vl_logic;
        A25             : in     vl_logic;
        A26             : in     vl_logic;
        A27             : in     vl_logic;
        A28             : in     vl_logic;
        A29             : in     vl_logic;
        A30             : in     vl_logic;
        A31             : in     vl_logic;
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        B4              : in     vl_logic;
        B5              : in     vl_logic;
        B6              : in     vl_logic;
        B7              : in     vl_logic;
        B8              : in     vl_logic;
        B9              : in     vl_logic;
        B10             : in     vl_logic;
        B11             : in     vl_logic;
        B12             : in     vl_logic;
        B13             : in     vl_logic;
        B14             : in     vl_logic;
        B15             : in     vl_logic;
        B16             : in     vl_logic;
        B17             : in     vl_logic;
        B18             : in     vl_logic;
        B19             : in     vl_logic;
        B20             : in     vl_logic;
        B21             : in     vl_logic;
        B22             : in     vl_logic;
        B23             : in     vl_logic;
        B24             : in     vl_logic;
        B25             : in     vl_logic;
        B26             : in     vl_logic;
        B27             : in     vl_logic;
        B28             : in     vl_logic;
        B29             : in     vl_logic;
        B30             : in     vl_logic;
        B31             : in     vl_logic;
        Cin             : in     vl_logic
    );
end Adder_32bit_nlogic;
