library verilog;
use verilog.vl_types.all;
entity TB_Adder_16bit is
end TB_Adder_16bit;
