library verilog;
use verilog.vl_types.all;
entity TB_Adder_32bit is
end TB_Adder_32bit;
