// Library - ECE555, Cell - INV_540_270, View - schematic
// LAST TIME SAVED: Oct 31 20:06:22 2011
// NETLIST TIME: Dec  1 16:12:42 2011
`timescale 1ns / 1ns 

module INV_540_270 ( OUT, IN );
output  OUT;

input  IN;


specify 
    specparam CDS_LIBNAME  = "ECE555";
    specparam CDS_CELLNAME = "INV_540_270";
    specparam CDS_VIEWNAME = "schematic";
endspecify

pmos P0 ( OUT, 1, IN);
nmos N0 ( OUT, 0, IN);

endmodule
